.MODEL 2N6755 NMOS( LEVEL=3 VTO=3.128 KP=21.14U PHI=600M GAMMA=0 TOX=100N 
+      UO=600 VMAX=0 DELTA=0 THETA=0 ETA=0 
+      L=2U W=1.1 RD=64.68M RS=120.7M RG=5.839 
+      RB=0 RDS=600K IS=44.14F N=1 PB=800M 
+      CBD=1.261N CBS=0 MJ=500M TT=370N CGSO=725.6P 
+      CGDO=310.6P CGBO=0 KF=0 AF=1 )


