.MODEL 1N5817 D( IS=1U N=537M BV=20 IBV=1M RS=55.6M 
+      CJO=210.8P VJ=0.35 M=1.442 FC=500M TT=1.67N 
+      EG=1.11 XTI=3 KF=0 AF=1 )

