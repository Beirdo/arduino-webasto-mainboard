.SUBCKT LMH6611  3 2 8 4 1
D17 9 0 DIN
D18 10 0 DIN
I14 0 9 0.1E-3
I15 0 10 0.1E-3
D19 11 0 DVN
D20 12 0 DVN
I16 0 11 0.1E-3
I17 0 12 0.1E-3
E15 13 2 11 12 2.6
G5 14 13 9 10 3E-4
E16 15 0 16 0 1
E17 17 0 18 0 1
E18 19 0 20 0 1
R56 15 21 1E6
R57 17 22 1E6
R58 19 23 1E6
R59 0 21 10
R60 0 22 10
R61 0 23 10
E19 24 25 23 0 1E-4
R62 26 20 1E3
R63 20 27 1E3
C15 15 21 1E-12
C16 17 22 1E-12
C17 19 23 1E-12
E20 28 24 22 0 -1
E21 29 28 21 0 2
R64 0 30 1E12
V52 30 0 1
G12 14 13 31 0 1.45E-14
R136 0 31 10E3
R137 0 31 10E3
R138 25 24 1E9
R139 24 28 1E9
R140 28 29 1E9
E54 27 0 14 0 1
E55 26 0 13 0 1
C23 14 13 0.25E-12
E57 25 3 32 0 2.25E-4
R146 25 3 1E9
R147 0 30 1E12
Q41 33 34 18 QLN
R148 34 35 1E3
R149 36 37 1E3
R150 38 16 1
R151 18 39 1
R153 40 41 5
R154 42 16 1
R155 18 43 1
D22 44 8 DD
D23 4 44 DD
E58 18 0 4 0 1
E59 16 0 8 0 1
R156 4 8 30E3
E60 45 18 16 18 0.5
D24 40 16 DD
D25 18 40 DD
R157 46 47 100
R158 48 49 100
G14 40 45 50 45 1E-3
R159 45 40 2E6
C24 41 51 3E-12
C25 44 0 1E-12
D26 49 33 DD
D27 52 47 DD
Q42 52 37 16 QLP
R160 44 53 1
R161 54 44 1
E61 55 45 56 57 1
R162 55 50 1E4
C26 50 45 0.025P
G15 58 45 40 45 -1E-3
G16 45 59 40 45 1E-3
G17 45 60 61 18 1E-3
G18 62 45 16 63 1E-3
D28 62 58 DD
D29 59 60 DD
R163 58 62 100E6
R164 60 59 100E6
R165 62 16 1E3
R166 18 60 1E3
R167 59 45 1E6
R168 60 45 1E6
R169 45 62 1E6
R170 45 58 1E6
G19 8 4 30 0 2.72E-3
R171 45 50 1E9
R172 46 16 1E9
R173 18 48 1E9
G20 63 61 30 0 0.25E-3
I22 8 4 0.5E-16
L2 44 1 3E-9
R175 44 1 1E3
R176 63 16 1E8
R177 18 61 1E8
R178 39 49 1E8
R179 38 47 1E8
R180 0 30 1E9
E99 16 36 8 38 4.8
E100 35 18 39 4 4.8
E124 51 0 44 0 1
R719 40 51 2E8
I30 0 64 1E-3
D46 64 0 DD
R778 0 64 10E6
V127 64 32 0.65
R779 0 32 10E6
Q52 53 47 38 QLP
Q53 54 49 39 QLN
Q54 61 61 43 QLN
Q55 63 63 42 QLP
E144 16 46 16 62 1
E145 48 18 60 18 1
Q56 65 14 66 QIN
Q57 67 13 68 QIN
Q58 57 69 65 QIN
Q59 56 70 67 QIN
Q60 69 69 16 QIP
Q61 14 69 16 QIP
Q62 70 70 16 QIP
Q63 13 70 16 QIP
R780 57 71 1200
R781 56 71 1200
R782 72 66 350
R783 72 68 350
Q64 72 73 74 QTN
I33 0 75 1E-3
D49 75 0 DD
R787 0 75 10E6
V130 75 76 1.2301
R788 0 76 10E6
E150 77 0 76 0 -1.75
R789 0 77 10E6
R790 78 77 10E6
M3 78 79 0 0 NEN L=2U W=1000U
G22 74 73 78 0 12E-6
V132 80 0 1
R791 80 79 1E6
M4 79 81 0 0 NEN L=2U W=100U
V133 81 0 1
C109 57 56 70F
V134 71 16 0.4
C110 0 14 2E-12
C111 13 0 2E-12
G23 8 0 53 44 1
G24 4 0 44 54 -1
G25 8 4 32 0 -2.4E-3
Q65 82 82 14 QIP
Q66 83 82 82 QIP
Q67 84 84 83 QIP
Q68 14 14 84 QIP
R792 13 83 50
V136 74 18 -0.9
J1 85 14 85 JNC
J2 85 13 85 JNC
J3 14 86 14 JNC
J4 13 86 13 JNC
V137 16 85 1.65
V138 86 18 0
I34 14 0 5.7E-6
I35 13 0 5.7E-6
.MODEL DD D
.MODEL QIN NPN BF=235 RB=900
.MODEL QIP PNP BF=235
.MODEL QTN NPN
.MODEL DVN D KF=2.5E-15
.MODEL DIN D KF=8E-15
.MODEL QLN NPN
.MODEL QLP PNP
.MODEL JNC NJF IS=1E-18
.MODEL NEN NMOS KP=200U VTO=0.5 IS=1E-18
.ENDS

