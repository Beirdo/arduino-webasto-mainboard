.MODEL 2N6804 PMOS( LEVEL=3 VTO=-1.695 KP=10.41U PHI=600M GAMMA=0 TOX=100N 
+      UO=300 VMAX=0 DELTA=0 THETA=0 ETA=0 
+      L=2U W=1.2 RD=66.52M RS=153M RG=4.931 
+      RB=0 RDS=444.4MEG IS=5.483P N=3 PB=800M 
+      CBD=1.291N CBS=0 MJ=500M TT=295N CGSO=1.783N 
+      CGDO=134.9P CGBO=0 KF=0 AF=1 )
